//============================================================================
//  Ultratank port to MiSTer
//  Copyright (c) 2020 Aitor Pelaez - NeuroRulez
//  EMU level .sv based on Alan Steremberg - alanswx work
//
//   
//============================================================================

module emu
(
	//Master input clock
	input         CLK_50M,

	//Async reset from top-level module.
	//Can be used as initial reset.
	input         RESET,

	//Must be passed to hps_io module
	inout  [45:0] HPS_BUS,

	//Base video clock. Usually equals to CLK_SYS.
	output        VGA_CLK,

	//Multiple resolutions are supported using different VGA_CE rates.
	//Must be based on CLK_VIDEO
	output        VGA_CE,

	output  [7:0] VGA_R,
	output  [7:0] VGA_G,
	output  [7:0] VGA_B,
	output        VGA_HS,
	output        VGA_VS,
	output        VGA_DE,    // = ~(VBlank | HBlank)
	output        VGA_F1,

	//Base video clock. Usually equals to CLK_SYS.
	output        HDMI_CLK,

	//Multiple resolutions are supported using different HDMI_CE rates.
	//Must be based on CLK_VIDEO
	output        HDMI_CE,

	output  [7:0] HDMI_R,
	output  [7:0] HDMI_G,
	output  [7:0] HDMI_B,
	output        HDMI_HS,
	output        HDMI_VS,
	output        HDMI_DE,   // = ~(VBlank | HBlank)
	output  [1:0] HDMI_SL,   // scanlines fx

	//Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
	output  [7:0] HDMI_ARX,
	output  [7:0] HDMI_ARY,

	output        LED_USER,  // 1 - ON, 0 - OFF.

	// b[1]: 0 - LED status is system status OR'd with b[0]
	//       1 - LED status is controled solely by b[0]
	// hint: supply 2'b00 to let the system control the LED.
	output  [1:0] LED_POWER,
	output  [1:0] LED_DISK,

	output [15:0] AUDIO_L,
	output [15:0] AUDIO_R,
	output        AUDIO_S,    // 1 - signed audio samples, 0 - unsigned

	// Open-drain User port.
	// 0 - D+/RX
	// 1 - D-/TX
	// 2..6 - USR2..USR6
	// Set USER_OUT to 1 to read from USER_IN.
	output        USER_OSD,	
	output        USER_MODE,
	input   [6:0] USER_IN,
	output  [6:0] USER_OUT
);

assign VGA_F1    = 0;

wire   JOY_CLK, JOY_LOAD;
wire   JOY_DATA  = USER_IN[5];
assign USER_OUT  = |status[31:30] ? {5'b11111,JOY_CLK,JOY_LOAD} : '1;
assign USER_MODE = |status[31:30] ;
assign USER_OSD  = joydb15_1[10] & joydb15_1[6];

assign LED_USER  = ioctl_download;
assign LED_DISK  = 2'b00;
assign LED_POWER = 2'b00;

assign HDMI_ARX = status[1] ? 8'd16 : 8'd4;
assign HDMI_ARY = status[1] ? 8'd9  : 8'd3;


`include "build_id.v"
localparam CONF_STR = {
	"A.ULTRATNK;;",
	"O1,Aspect Ratio,Original,Wide;",
	"O35,Scandoubler Fx,None,HQ2x,CRT 25%,CRT 50%,CRT 75%;",  
	"OUV,Serial SNAC DB15,Off,1 Player,2 Players;",	
	"-;",
	"O89,Extended Play,none,25pts,50pts,75pts;",
	"OAB,Game time,150 Sec,120 Sec,90 Sec,60 Sec;",
	"OC,Color,Off,On;",
	"OD,Test,Off,On;",
	"OE,Invisible tanks,Off,On;",
	"OF,Rebounding shells,Off,On;",
	"OG,Barriers,On,Off;",
	"-;",
	"R0,Reset;",
	"J1,Fire,Start 1P,Start 2P,Coin;",
	"V,v",`BUILD_DATE
};



wire [31:0] status;
wire  [1:0] buttons;
wire        ioctl_download;
wire        ioctl_wr;
wire [24:0] ioctl_addr;
wire [7:0] ioctl_data;

wire        forced_scandoubler;
wire [21:0] gamma_bus;
wire [10:0] ps2_key;

wire [15:0] joy1_USB, joy2_USB;

wire [31:0] joy1 = |status[31:30] ? {joydb15_1[11],joydb15_1[9],joydb15_1[10],joydb15_1[4:0]} : joy1_USB;
wire [31:0] joy2 =  status[31]    ? {joydb15_2[11],joydb15_2[10],joydb15_2[9],joydb15_2[4:0]} : status[30] ? joy1_USB : joy2_USB;

//----BA 9876543210
//----LS FEDCBAUDLR
reg [15:0] joydb15_1,joydb15_2;
joy_db15 joy_db15
(
  .clk       ( CLK_50M   ), //48MHz
  .JOY_CLK   ( JOY_CLK   ),
  .JOY_DATA  ( JOY_DATA  ),
  .JOY_LOAD  ( JOY_LOAD  ),
  .joystick1 ( joydb15_1 ),
  .joystick2 ( joydb15_2 )	  
);


hps_io #(.STRLEN(($size(CONF_STR)>>3) )) hps_io
(
	.clk_sys(clk_sys),
	.HPS_BUS(HPS_BUS),

	.conf_str(CONF_STR),
	
	.buttons(buttons),
	.status(status),
	.forced_scandoubler(forced_scandoubler),
	.gamma_bus(gamma_bus),


	.ioctl_download(ioctl_download),
	.ioctl_wr(ioctl_wr),
	.ioctl_addr(ioctl_addr),
	.ioctl_dout(ioctl_data),
	
	.joy_raw(joydb15_1[5:0]),
	.joystick_0(joy1_USB),
	.joystick_1(joy2_USB),
	.ps2_key(ps2_key)
);



wire       pressed = ps2_key[9];
wire [8:0] code    = ps2_key[8:0];
always @(posedge clk_sys) begin
	reg old_state;
	old_state <= ps2_key[10];
	
	if(old_state != ps2_key[10]) begin
		casex(code)
			'hX75: btn_up          <= pressed; // up
			'hX72: btn_down        <= pressed; // down
			'hX6B: btn_left        <= pressed; // left
			'hX74: btn_right       <= pressed; // right
			'h014: btn_fire        <= pressed; // ctrl			

			'h005: btn_one_player  <= pressed; // F1
			'h006: btn_two_players <= pressed; // F2
			'h004: btn_coin        <= pressed; // F3
			
			// JPAC/IPAC/MAME Style Codes
			'h016: btn_start_1     <= pressed; // 1
			'h01E: btn_start_2     <= pressed; // 2
			'h02E: btn_coin_1      <= pressed; // 5
			'h036: btn_coin_2      <= pressed; // 6

			'h02D: btn_up_2        <= pressed; // R
			'h02B: btn_down_2      <= pressed; // F
			'h023: btn_left_2      <= pressed; // D
			'h034: btn_right_2     <= pressed; // G
			'h01C: btn_fire_2      <= pressed; // A
		endcase
	end
end

reg btn_up    = 0;
reg btn_down  = 0;
reg btn_right = 0;
reg btn_left  = 0;
reg btn_fire  = 0;

reg btn_one_player  = 0;
reg btn_two_players = 0;

reg btn_start_1=0;
reg btn_start_2=0;
reg btn_coin  = 0;
reg btn_coin_1=0;
reg btn_coin_2=0;
reg btn_up_2=0;
reg btn_down_2=0;
reg btn_left_2=0;
reg btn_right_2=0;
reg btn_fire_2=0;

wire m_fire     = btn_fire    | joy1[4];
wire m_fire_2   = btn_fire_2  | joy2[4];
wire m_start    = btn_start_1 | joy1[5] | joy2[5];
wire m_start_2  = btn_start_2 | joy1[6] | joy2[6];
wire m_coin     = btn_coin    | joy1[7] | joy2[7] | btn_coin_1 | btn_coin_2;

wire m_up      = btn_up      | joy1[3];
wire m_down    = btn_down    | joy1[2];
wire m_left    = btn_left    | joy1[1];
wire m_right   = btn_right   | joy1[0];
wire m_up_2    = btn_up_2    | joy2[3];
wire m_down_2  = btn_down_2  | joy2[2];
wire m_left_2  = btn_left_2  | joy2[1];
wire m_right_2 = btn_right_2 | joy2[0];


wire compositesync;
wire [5:0] video_r,video_g,video_b;

tld_test_placa_mister tld_test_placa_mister(
	.clk7(clk_7),
	//.Reset_n(~(RESET | status[0]  | buttons[1] | ioctl_download)),
	.BTN_USER(~btn_one_player),

	.r_to_vga(r),
	.g_to_vga(g),
	.b_to_vga(b),

	.hsync_to_vga(hs),
	.vsync_to_vga(vs),
	.hblank_to_vga(hblank),
	.vblank_to_vga(vblank),
	.csync_to_vga(compositesync),
	
	.joy1(joydb15_1),
	.joy2(joydb15_2),
	
	.CLK_VIDEO(CLK_VIDEO_2)
	);
			
wire [6:0] audio1;
wire [6:0] audio2;
wire [1:0] video;
wire [3:0] videor;
///////////////////////////////////////////////////
wire clk_14,clk_7,CLK_VIDEO_2;
wire clk_sys,locked;

assign AUDIO_L={audio1,1'b0,8'b00000000};
assign AUDIO_R={audio2,1'b0,8'b00000000};
assign AUDIO_S = 0;

wire hblank, vblank;
wire hs, vs;
wire [5:0] r,g,b;

reg ce_pix;
always @(posedge clk_14) begin
        reg old_clk;

        old_clk <= CLK_VIDEO_2;
        ce_pix <= old_clk & ~CLK_VIDEO_2;
end

arcade_video #(320,9) arcade_video
(
        .*,

        .clk_video(clk_14),

        .RGB_in({r,g,b}),
        .HBlank(hblank),
        .VBlank(vblank),
        .HSync(hs),
        .VSync(vs),

        .fx(status[5:3]),
		  .rotate_ccw(0),
	     .no_rotate(1)		  
);

pll pll (
	.refclk ( CLK_50M   ),
	.rst(0),
	.locked 		( locked    ),        // PLL is running stable
	.outclk_0	( clk_14	),        // 24 MHz
	.outclk_1	( clk_7  	)        // 7 MHz
	 );

assign clk_sys=clk_14;

endmodule
